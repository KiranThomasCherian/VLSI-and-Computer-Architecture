magic
tech scmos
timestamp 1597230813
<< nwell >>
rect -12 17 35 31
<< polysilicon >>
rect 1 29 4 35
rect 18 29 21 35
rect 1 -3 4 19
rect 18 -3 21 19
rect 1 -17 4 -13
rect 18 -17 21 -13
<< ndiffusion >>
rect -10 -6 1 -3
rect -10 -12 -7 -6
rect -1 -12 1 -6
rect -10 -13 1 -12
rect 4 -6 18 -3
rect 4 -12 8 -6
rect 14 -12 18 -6
rect 4 -13 18 -12
rect 21 -6 33 -3
rect 21 -12 24 -6
rect 30 -12 33 -6
rect 21 -13 33 -12
<< pdiffusion >>
rect -10 28 1 29
rect -10 22 -7 28
rect 0 22 1 28
rect -10 19 1 22
rect 4 19 18 29
rect 21 26 33 29
rect 21 20 22 26
rect 28 20 33 26
rect 21 19 33 20
<< metal1 >>
rect -7 38 -6 44
rect 0 38 7 44
rect 13 38 20 44
rect 26 38 28 44
rect -7 37 28 38
rect -7 28 0 37
rect 22 13 28 20
rect 8 8 28 13
rect 8 -6 15 8
rect 14 -12 15 -6
rect 24 -6 30 -5
rect -7 -19 -1 -12
rect 24 -19 30 -12
rect -1 -24 4 -19
rect 10 -24 14 -19
rect 20 -24 24 -19
<< ntransistor >>
rect 1 -13 4 -3
rect 18 -13 21 -3
<< ptransistor >>
rect 1 19 4 29
rect 18 19 21 29
<< ndcontact >>
rect -7 -12 -1 -6
rect 8 -12 14 -6
rect 24 -12 30 -6
<< pdcontact >>
rect -7 22 0 28
rect 22 20 28 26
<< psubstratepcontact >>
rect -7 -24 -1 -19
rect 4 -24 10 -19
rect 14 -24 20 -19
rect 24 -24 30 -19
<< nsubstratencontact >>
rect -6 38 0 44
rect 7 38 13 44
rect 20 38 26 44
<< labels >>
rlabel polysilicon 2 3 2 3 1 A
rlabel polysilicon 20 3 20 3 1 B
rlabel metal1 26 11 26 11 1 Y
rlabel metal1 4 41 4 41 5 vdd
rlabel metal1 1 -22 1 -22 1 gnd
<< end >>
