//`include "adder32_a.v"
`include "Myfinal_32cla.v"
module cla_testbench;
reg [31:0] a, b;
reg cin;
wire [31:0] sum;
wire cout;

thirtytwo_bit_Recursive_Carry_Adder adder(sum[31:0],cout,a[31:0],b[31:0]);
initial
begin
  $display("	a +	b	=	sum 	,	carryout");
end
    
initial
begin
     a='b11111111111111111111111111111111; b='b11111111111111111111111111111111;
  #30 a='b00000000000000000000000000000000; b='b11111111111111111111111111111111;
  #30 a='b10101010101010101010101010101010; b='b01010101010101010101010101010101;
  #30 a='b11001100110011001100110011001100; b='b11000000000001100000000000111101;
  #30 a='b11001100110011001100110011001100; b='b00000000000000000000111111111111; 
  #30 a='b10000000000000000000000000000001; b='b10000000000000000000000000000111;
  #30 a='b0000; b='b00111;

end

initial
begin
  $monitor(" %b + %b = %b cout= %b ", a[31:0],b[31:0],sum[31:0],cout);
end
endmodule
