`include "Float_multiply.v"
module tb;

reg [31:0] a,b;
wire[31:0] out;
reg clk;
fmultiplier m1(out,a,b,clk);

initial 
begin
		clk = 0;
		forever begin
			#5 clk = ~clk;
		end
end
initial 
begin
	 a=32'b01000011010010001100000000000000; b=32'b01111111100000000000000000000000; //infinity
    #10 a=32'b01000001000111000000000000000000; b=32'b00111111000100000000000000000000;	 //9.75 and 0.5625
	#10 a=32'b01000001010010000000000000000000; b=32'b11000000101100100000000000000000;  //12.5 and -5.5625		-69.53125 

  #10 b = 32'b01111111100000000000000000000001; //nan
   #10     a=32'b00000000000000000000000000000000; b=32'b01000000101000000000000000000000;


    #500 $finish;
end
initial
    $monitor($time," a = %b * b = %b ; out = %b ;",a,b,out);

endmodule
